* Created by KLayout

* cell nand
* pin B
* pin A
* pin Z
* pin VSS
* pin VDD
.SUBCKT nand 1 3 4 5 6
* net 1 B
* net 3 A
* net 4 Z
* net 5 VSS
* net 6 VDD
* device instance $1 r0 *1 1067,-222.5 NMOS
M$1 43 47 45 43 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $2 r0 *1 1067,-382.5 NMOS
M$2 44 48 46 44 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $3 r0 *1 907,-222.5 NMOS
M$3 16 22 34 16 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $4 r0 *1 907,-382.5 NMOS
M$4 19 37 13 19 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $5 r0 *1 1067,-862.5 NMOS
M$5 49 53 51 49 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $6 r0 *1 1067,-1022.5 NMOS
M$6 50 54 52 50 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $7 r0 *1 907,-862.5 NMOS
M$7 17 23 35 17 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $8 r0 *1 907,-1022.5 NMOS
M$8 20 38 14 20 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $9 r0 *1 427,-222.5 NMOS
M$9 55 59 57 55 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $10 r0 *1 427,-382.5 NMOS
M$10 56 60 58 56 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $11 r0 *1 267,-222.5 NMOS
M$11 4 3 2 4 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $12 r0 *1 267,-382.5 NMOS
M$12 4 1 5 4 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $13 r0 *1 427,-862.5 NMOS
M$13 61 65 63 61 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $14 r0 *1 427,-1022.5 NMOS
M$14 62 66 64 62 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $15 r0 *1 267,-862.5 NMOS
M$15 18 24 36 18 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $16 r0 *1 267,-1022.5 NMOS
M$16 21 39 15 21 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $17 r0 *1 1070,114 PMOS
M$17 69 71 67 69 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $18 r0 *1 1070,-46 PMOS
M$18 70 72 68 70 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $19 r0 *1 910,114 PMOS
M$19 28 40 10 28 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $20 r0 *1 910,-46 PMOS
M$20 31 25 7 31 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $21 r0 *1 1070,-526 PMOS
M$21 75 77 73 75 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $22 r0 *1 1070,-686 PMOS
M$22 76 78 74 76 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $23 r0 *1 910,-526 PMOS
M$23 29 41 11 29 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $24 r0 *1 910,-686 PMOS
M$24 32 26 8 32 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $25 r0 *1 430,114 PMOS
M$25 81 83 79 81 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $26 r0 *1 430,-46 PMOS
M$26 82 84 80 82 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $27 r0 *1 270,114 PMOS
M$27 2 1 6 2 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $28 r0 *1 270,-46 PMOS
M$28 2 3 6 2 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $29 r0 *1 430,-526 PMOS
M$29 87 89 85 87 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $30 r0 *1 430,-686 PMOS
M$30 88 90 86 88 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $31 r0 *1 270,-526 PMOS
M$31 30 42 12 30 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $32 r0 *1 270,-686 PMOS
M$32 33 27 9 33 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
.ENDS nand
