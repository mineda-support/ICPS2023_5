* Created by KLayout

* cell nand
.SUBCKT nand
* device instance $1 r0 *1 1067,-222.5 NMOS
M$1 45 47 43 43 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $2 r0 *1 1067,-382.5 NMOS
M$2 46 48 44 44 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $3 r0 *1 907,-222.5 NMOS
M$3 34 22 16 16 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $4 r0 *1 907,-382.5 NMOS
M$4 13 37 19 19 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $5 r0 *1 1067,-862.5 NMOS
M$5 51 53 49 49 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $6 r0 *1 1067,-1022.5 NMOS
M$6 52 54 50 50 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $7 r0 *1 907,-862.5 NMOS
M$7 35 23 17 17 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $8 r0 *1 907,-1022.5 NMOS
M$8 14 38 20 20 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $9 r0 *1 427,-222.5 NMOS
M$9 57 59 55 55 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $10 r0 *1 427,-382.5 NMOS
M$10 58 60 56 56 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $11 r0 *1 267,-222.5 NMOS
M$11 2 3 4 4 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $12 r0 *1 267,-382.5 NMOS
M$12 5 1 4 4 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $13 r0 *1 427,-862.5 NMOS
M$13 63 65 61 61 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $14 r0 *1 427,-1022.5 NMOS
M$14 64 66 62 62 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $15 r0 *1 267,-862.5 NMOS
M$15 36 24 18 18 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $16 r0 *1 267,-1022.5 NMOS
M$16 15 39 21 21 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $17 r0 *1 1070,114 PMOS
M$17 67 71 69 69 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $18 r0 *1 1070,-46 PMOS
M$18 68 72 70 70 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $19 r0 *1 910,114 PMOS
M$19 10 40 28 28 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $20 r0 *1 910,-46 PMOS
M$20 7 25 31 31 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $21 r0 *1 1070,-526 PMOS
M$21 73 77 75 75 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $22 r0 *1 1070,-686 PMOS
M$22 74 78 76 76 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $23 r0 *1 910,-526 PMOS
M$23 11 41 29 29 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $24 r0 *1 910,-686 PMOS
M$24 8 26 32 32 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $25 r0 *1 430,114 PMOS
M$25 79 83 81 81 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $26 r0 *1 430,-46 PMOS
M$26 80 84 82 82 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $27 r0 *1 270,114 PMOS
M$27 6 1 2 2 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $28 r0 *1 270,-46 PMOS
M$28 6 3 2 2 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $29 r0 *1 430,-526 PMOS
M$29 85 89 87 87 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $30 r0 *1 430,-686 PMOS
M$30 86 90 88 88 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $31 r0 *1 270,-526 PMOS
M$31 12 42 30 30 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
* device instance $32 r0 *1 270,-686 PMOS
M$32 9 27 33 33 PMOS L=10U W=40U AS=760P AD=760P PS=118U PD=118U
.ENDS nand
